module tb;
wire k;
task3 u0(.k(k));
initial begin
u0.display();
end
endmodule
