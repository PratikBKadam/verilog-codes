module fabehave(a,b,c0,s,c);
input a,b,c0;
output reg s,c;
always @(*)
begin
if(c0)
begin
if(a)
begin
if(b)
begin
s=1'b1;
c=1'b1;
end
else
begin
s=1'b0;
c=1'b1;
end
end
else
begin
if(b)
begin
s=1'b0;
c=1'b1;
end
else
begin
s=1'b1;
c=1'b0;
end
end
end
else
begin
if(a)
begin
if(b)
begin
s=1'b0;
c=1'b1;
end
else
begin
s=1'b1;
c=1'b0;
end
end
else
begin
if(b)
begin
s=1'b1;
c=1'b0;
end
else
begin
s=1'b0;
c=1'b0;
end
end
end
end
endmodule
