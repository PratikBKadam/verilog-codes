module task3(output k);
task display;
begin
$display("-");
end
endtask
display();

assign k=0;
endmodule
